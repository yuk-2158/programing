timescale 1ns/1ps
//Module Name: full_adder_by_elements

module full_adder_by_elements(
  input wire x2, x1, x0,
  output wire[1:0] y
);
  assign y[1] =  ;
  assign y[0] =   ;
endmodule
  
